module gpu_cache_L1(
	input wire clk,
	output wire out
	);

endmodule